module ast

pub interface Stmt {
	stmt()
}

pub interface Expr {
	expr()
}